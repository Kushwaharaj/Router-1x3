module router_synchronizer(clock,resetn,detect_add,write_enb_reg,read_enb_0,read_enb_1,read_enb_2,data_in,
full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb,vld_out_0,vld_out_1,vld_out_2,soft_reset_0,soft_reset_1,soft_reset_2,fifo_full);
input clock,resetn,detect_add,write_enb_reg,read_enb_0,read_enb_1,read_enb_2,full_0,full_1,full_2,empty_0,empty_1,empty_2;
input [1:0] data_in;
output reg [2:0] write_enb;
output reg soft_reset_0,soft_reset_1,soft_reset_2,fifo_full;
output vld_out_0,vld_out_1,vld_out_2;
reg [1:0] temp;
reg [4:0] count_0,count_1,count_2;
//generating valid out signal if the FIFO is empty and it can accept data
assign vld_out_0 = ~empty_0;
assign vld_out_1 = ~empty_1;
assign vld_out_2 = ~empty_2;

//fetching the address and storing in a temporary variable
always@(posedge clock)
begin
if(!resetn)
temp<=0;
else if(detect_add)
temp<=data_in;
end

//Logic for fifo_full signal based on which of the fifo is full
always@(*)
begin
case(temp)
2'b00:fifo_full=full_0;
2'b01:fifo_full=full_1;
2'b10:fifo_full=full_2;
default:fifo_full=1'b0;
endcase
end

//if write_enb_reg is high then generate write enable signal(one hot encoding) for that FIFO
always@(*)
begin
if(write_enb_reg)
begin
case(temp)
2'b00:write_enb=3'b001;
2'b01:write_enb=3'b010;
2'b10:write_enb=3'b100;
default:write_enb=3'b000;
endcase
end
else
write_enb=3'b000;
end

//once read_enable is asserted,reset the counter to 0
always@(posedge clock)
 begin
  if(!resetn)
    count_0<=5'b0;

  else if(vld_out_0)
    begin
      if(!read_enb_0)
        begin
          if(count_0==29)
            begin
              soft_reset_0<=1'b1;
              count_0<=5'b0;
            end
          else
            begin
              count_0<=count_0+5'b1;
              soft_reset_0<=1'b0;
            end
        end
      else count_0<=5'b0;
    end
  else count_0<=5'b0;
end

always@(posedge clock)
begin
if(!resetn)
count_1<=5'b0;

else if(vld_out_1)
begin
if(!read_enb_1)
begin
if(count_1==29)
begin
soft_reset_1<=1'b1;
count_1<=5'b0;
end
else
begin
count_1<=count_1+5'b1;
soft_reset_1<=1'b0;
end
end
else count_1<=5'b0;
end
else count_1<=5'b0;
end

always@(posedge clock)
begin
if(!resetn)
count_2<=5'b0;

else if(vld_out_2)
begin
if(!read_enb_2)
begin
if(count_2==29)
begin
soft_reset_2<=1'b1;
count_2<=5'b0;
end
else
begin
count_2<=count_2+5'b1;
soft_reset_2<=1'b0;
end
end
else count_2<=5'b0;
end
else count_2<=5'b0;
end
endmodule
